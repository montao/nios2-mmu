// qsys.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module qsys (
		input  wire        clk_clk,                      //                      clk.clk
		input  wire        reset_reset_n,                //                    reset.reset_n
		output wire [12:0] sdram_wire_addr,              //               sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                //                         .ba
		output wire        sdram_wire_cas_n,             //                         .cas_n
		output wire        sdram_wire_cke,               //                         .cke
		output wire        sdram_wire_cs_n,              //                         .cs_n
		inout  wire [31:0] sdram_wire_dq,                //                         .dq
		output wire [3:0]  sdram_wire_dqm,               //                         .dqm
		output wire        sdram_wire_ras_n,             //                         .ras_n
		output wire        sdram_wire_we_n,              //                         .we_n
		input  wire        uart_external_connection_rxd, // uart_external_connection.rxd
		output wire        uart_external_connection_txd  //                         .txd
	);

	wire  [31:0] cpu_data_master_readdata;                             // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                          // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                          // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                              // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                           // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                 // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                        // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                            // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                      // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                   // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                       // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                          // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                 // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;       // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;    // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;        // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;           // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;          // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_mmu_s1_chipselect;              // mm_interconnect_0:ram_mmu_s1_chipselect -> ram_mmu:chipselect
	wire  [31:0] mm_interconnect_0_ram_mmu_s1_readdata;                // ram_mmu:readdata -> mm_interconnect_0:ram_mmu_s1_readdata
	wire   [7:0] mm_interconnect_0_ram_mmu_s1_address;                 // mm_interconnect_0:ram_mmu_s1_address -> ram_mmu:address
	wire   [3:0] mm_interconnect_0_ram_mmu_s1_byteenable;              // mm_interconnect_0:ram_mmu_s1_byteenable -> ram_mmu:byteenable
	wire         mm_interconnect_0_ram_mmu_s1_write;                   // mm_interconnect_0:ram_mmu_s1_write -> ram_mmu:write
	wire  [31:0] mm_interconnect_0_ram_mmu_s1_writedata;               // mm_interconnect_0:ram_mmu_s1_writedata -> ram_mmu:writedata
	wire         mm_interconnect_0_ram_mmu_s1_clken;                   // mm_interconnect_0:ram_mmu_s1_clken -> ram_mmu:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                  // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;               // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                   // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                      // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;             // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                     // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                 // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_s1_chipselect;                // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                  // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                   // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                     // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                 // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                 // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                   // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                    // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                       // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;              // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                      // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                  // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_ram_mmu_s2_chipselect;              // mm_interconnect_0:ram_mmu_s2_chipselect -> ram_mmu:chipselect2
	wire  [31:0] mm_interconnect_0_ram_mmu_s2_readdata;                // ram_mmu:readdata2 -> mm_interconnect_0:ram_mmu_s2_readdata
	wire   [7:0] mm_interconnect_0_ram_mmu_s2_address;                 // mm_interconnect_0:ram_mmu_s2_address -> ram_mmu:address2
	wire   [3:0] mm_interconnect_0_ram_mmu_s2_byteenable;              // mm_interconnect_0:ram_mmu_s2_byteenable -> ram_mmu:byteenable2
	wire         mm_interconnect_0_ram_mmu_s2_write;                   // mm_interconnect_0:ram_mmu_s2_write -> ram_mmu:write2
	wire  [31:0] mm_interconnect_0_ram_mmu_s2_writedata;               // mm_interconnect_0:ram_mmu_s2_writedata -> ram_mmu:writedata2
	wire         mm_interconnect_0_ram_mmu_s2_clken;                   // mm_interconnect_0:ram_mmu_s2_clken -> ram_mmu:clken2
	wire         irq_mapper_receiver0_irq;                             // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                             // uart:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                          // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, jtag:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, ram_mmu:reset, ram_mmu:reset2, rst_translator:in_reset, sdram:reset_n, timer:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [cpu:reset_req, ram_mmu:reset_req, ram_mmu:reset_req2, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                        // cpu:debug_reset_request -> rst_controller:reset_in1

	qsys_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	qsys_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	qsys_ram_mmu ram_mmu (
		.clk         (clk_clk),                                 //   clk1.clk
		.address     (mm_interconnect_0_ram_mmu_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_ram_mmu_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_ram_mmu_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_ram_mmu_s1_write),      //       .write
		.readdata    (mm_interconnect_0_ram_mmu_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_ram_mmu_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_ram_mmu_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.address2    (mm_interconnect_0_ram_mmu_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_ram_mmu_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_ram_mmu_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_ram_mmu_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_ram_mmu_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_ram_mmu_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_ram_mmu_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                 //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),          // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze      (1'b0)                                     // (terminated)
	);

	qsys_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	qsys_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	qsys_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_external_connection_rxd),            // external_connection.export
		.txd           (uart_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                        (clk_clk),                                              //                      clk_50_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address               (cpu_data_master_address),                              //                 cpu_data_master.address
		.cpu_data_master_waitrequest           (cpu_data_master_waitrequest),                          //                                .waitrequest
		.cpu_data_master_byteenable            (cpu_data_master_byteenable),                           //                                .byteenable
		.cpu_data_master_read                  (cpu_data_master_read),                                 //                                .read
		.cpu_data_master_readdata              (cpu_data_master_readdata),                             //                                .readdata
		.cpu_data_master_readdatavalid         (cpu_data_master_readdatavalid),                        //                                .readdatavalid
		.cpu_data_master_write                 (cpu_data_master_write),                                //                                .write
		.cpu_data_master_writedata             (cpu_data_master_writedata),                            //                                .writedata
		.cpu_data_master_debugaccess           (cpu_data_master_debugaccess),                          //                                .debugaccess
		.cpu_instruction_master_address        (cpu_instruction_master_address),                       //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                   //                                .waitrequest
		.cpu_instruction_master_read           (cpu_instruction_master_read),                          //                                .read
		.cpu_instruction_master_readdata       (cpu_instruction_master_readdata),                      //                                .readdata
		.cpu_instruction_master_readdatavalid  (cpu_instruction_master_readdatavalid),                 //                                .readdatavalid
		.cpu_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),        //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),          //                                .write
		.cpu_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),           //                                .read
		.cpu_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),       //                                .readdata
		.cpu_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),      //                                .writedata
		.cpu_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),     //                                .byteenable
		.cpu_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),    //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),    //                                .debugaccess
		.jtag_avalon_jtag_slave_address        (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //          jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write          (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                .write
		.jtag_avalon_jtag_slave_read           (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                .read
		.jtag_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                .chipselect
		.ram_mmu_s1_address                    (mm_interconnect_0_ram_mmu_s1_address),                 //                      ram_mmu_s1.address
		.ram_mmu_s1_write                      (mm_interconnect_0_ram_mmu_s1_write),                   //                                .write
		.ram_mmu_s1_readdata                   (mm_interconnect_0_ram_mmu_s1_readdata),                //                                .readdata
		.ram_mmu_s1_writedata                  (mm_interconnect_0_ram_mmu_s1_writedata),               //                                .writedata
		.ram_mmu_s1_byteenable                 (mm_interconnect_0_ram_mmu_s1_byteenable),              //                                .byteenable
		.ram_mmu_s1_chipselect                 (mm_interconnect_0_ram_mmu_s1_chipselect),              //                                .chipselect
		.ram_mmu_s1_clken                      (mm_interconnect_0_ram_mmu_s1_clken),                   //                                .clken
		.ram_mmu_s2_address                    (mm_interconnect_0_ram_mmu_s2_address),                 //                      ram_mmu_s2.address
		.ram_mmu_s2_write                      (mm_interconnect_0_ram_mmu_s2_write),                   //                                .write
		.ram_mmu_s2_readdata                   (mm_interconnect_0_ram_mmu_s2_readdata),                //                                .readdata
		.ram_mmu_s2_writedata                  (mm_interconnect_0_ram_mmu_s2_writedata),               //                                .writedata
		.ram_mmu_s2_byteenable                 (mm_interconnect_0_ram_mmu_s2_byteenable),              //                                .byteenable
		.ram_mmu_s2_chipselect                 (mm_interconnect_0_ram_mmu_s2_chipselect),              //                                .chipselect
		.ram_mmu_s2_clken                      (mm_interconnect_0_ram_mmu_s2_clken),                   //                                .clken
		.sdram_s1_address                      (mm_interconnect_0_sdram_s1_address),                   //                        sdram_s1.address
		.sdram_s1_write                        (mm_interconnect_0_sdram_s1_write),                     //                                .write
		.sdram_s1_read                         (mm_interconnect_0_sdram_s1_read),                      //                                .read
		.sdram_s1_readdata                     (mm_interconnect_0_sdram_s1_readdata),                  //                                .readdata
		.sdram_s1_writedata                    (mm_interconnect_0_sdram_s1_writedata),                 //                                .writedata
		.sdram_s1_byteenable                   (mm_interconnect_0_sdram_s1_byteenable),                //                                .byteenable
		.sdram_s1_readdatavalid                (mm_interconnect_0_sdram_s1_readdatavalid),             //                                .readdatavalid
		.sdram_s1_waitrequest                  (mm_interconnect_0_sdram_s1_waitrequest),               //                                .waitrequest
		.sdram_s1_chipselect                   (mm_interconnect_0_sdram_s1_chipselect),                //                                .chipselect
		.timer_s1_address                      (mm_interconnect_0_timer_s1_address),                   //                        timer_s1.address
		.timer_s1_write                        (mm_interconnect_0_timer_s1_write),                     //                                .write
		.timer_s1_readdata                     (mm_interconnect_0_timer_s1_readdata),                  //                                .readdata
		.timer_s1_writedata                    (mm_interconnect_0_timer_s1_writedata),                 //                                .writedata
		.timer_s1_chipselect                   (mm_interconnect_0_timer_s1_chipselect),                //                                .chipselect
		.uart_s1_address                       (mm_interconnect_0_uart_s1_address),                    //                         uart_s1.address
		.uart_s1_write                         (mm_interconnect_0_uart_s1_write),                      //                                .write
		.uart_s1_read                          (mm_interconnect_0_uart_s1_read),                       //                                .read
		.uart_s1_readdata                      (mm_interconnect_0_uart_s1_readdata),                   //                                .readdata
		.uart_s1_writedata                     (mm_interconnect_0_uart_s1_writedata),                  //                                .writedata
		.uart_s1_begintransfer                 (mm_interconnect_0_uart_s1_begintransfer),              //                                .begintransfer
		.uart_s1_chipselect                    (mm_interconnect_0_uart_s1_chipselect)                  //                                .chipselect
	);

	qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
